// GAME CONSTANTS
parameter MAX_X = 127;
parameter MIN_X = 0;
parameter MAX_Y = 95;
parameter MIN_Y = 0;
parameter LEFT = 0;
parameter RIGHT = 1;

// PLAYER STATES
parameter NUM_STATES = 8;

parameter DEFAULT_STATE = 0;
parameter JUMP_STATE = 1;
parameter CROUCH_STATE = 2;
parameter MELEE_STATE_LEFT = 3;
parameter RANGED_STATE = 4;
parameter HIT_STATE = 5;
parameter MELEE_STATE_RIGHT = 6;

// FIREBALL STATES
parameter FIREBALL_DISABLED = 0;
parameter FIREBALL_ENABLED = 1;
parameter FIREBALL_EXPLOSION = 2;

// Y-LEVELS
parameter GROUND_LEVEL = 70;
parameter JUMP_LEVEL = 10;

// COLORS
parameter SKY_BLUE = 8'd50;
parameter LIGHT_GREEN = 8'd20;
parameter WHITE = 8'd255;
parameter BLACK = 8'd0;
parameter RED = 8'd224;
parameter GREEN = 8'd28;
parameter BLUE = 8'd3;
parameter ORANGE = 8'd236;

// SPRITES
parameter SPRITE_HEIGHT = 4;
parameter SPRITE_WIDTH = 3;

const logic [0:NUM_STATES-1][0:SPRITE_HEIGHT-1][0:SPRITE_WIDTH-1][7:0] SPRITE = {

    // DEFAULT STATE:
    {   SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , BLACK     , BLACK,
        SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , SKY_BLUE  , BLACK         },

    // JUMP STATE:
    {   SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , BLACK     , BLACK,
        BLACK       , BLACK     , BLACK,
        BLACK       , SKY_BLUE  , BLACK         },

    // CROUCH STATE:
    {   SKY_BLUE    , SKY_BLUE  , SKY_BLUE,
        SKY_BLUE    , SKY_BLUE  , SKY_BLUE,
        BLACK       , BLACK     , BLACK,
        BLACK       , BLACK     , BLACK         },

    // MELEE STATE LEFT:
    {   SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , BLACK     , SKY_BLUE,
        SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , SKY_BLUE  , BLACK         },

    // RANGED STATE:
    {   SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , BLACK     , BLACK,
        SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , SKY_BLUE  , BLACK         },

    // HIT STATE:
    {   SKY_BLUE    , RED       , SKY_BLUE,
        RED         , RED       , RED,
        SKY_BLUE    , RED       , SKY_BLUE,
        RED         , SKY_BLUE  , RED           },

    // MELEEE STATE RIGHT:
    {   SKY_BLUE    , BLACK     , SKY_BLUE,
        SKY_BLUE    , BLACK     , BLACK,
        SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , SKY_BLUE  , BLACK         },

    // 
    {   SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , BLACK     , BLACK,
        SKY_BLUE    , BLACK     , SKY_BLUE,
        BLACK       , SKY_BLUE  , BLACK         }

};


const logic [0:17][0:32] GAME_OVER_BITMAP = {
    33'b000000000000000000000000000000000,
    33'b000111110001110001100011011111110,
    33'b001100000011011001110111011000000,
    33'b011000000110001101111111011000000,
    33'b011001110110001101111111011111100,
    33'b011000110111111101101011011000000,
    33'b001100110110001101100011011000000,
    33'b000111110110001101100011011111110,
    33'b000000000000000000000000000000000,
    33'b000000000000000000000000000000000,
    33'b001111100110001101111111011111100,
    33'b011000110110001101100000011000110,
    33'b011000110110001101100000011000110,
    33'b011000110111011101111110011001110,
    33'b011000110011111001100000011111000,
    33'b011000110001110001100000011011100,
    33'b001111100000100001111111011001110,
    33'b000000000000000000000000000000000
};

const logic [0:8][0:71] PLAYER_BLANK_WINS_BITMAP = {    
    //  PPPPP LL AAAAA YYYYY EEEE RRRR      1or2      WWWWWWW II NNNNN SSSS   !!
    72'b000000000000000000000000000000000000000000000000000000000000000000000011,
    72'b000000110000000000000000000000000000000000000000000000110000000000000011,
    72'b000000110000000000000000000000000000000000000000000000000000000000000011,
    72'b111110110111100100110111101111000000000000000011000110110111100111100011,
    72'b110010110100110100110111101101000000000000000011010110110110010110000011,
    72'b110010110100110100110100001100000000000000000011111110110110010001100000,
    72'b111110110111110111110111101100000000000000000001101100110110010111100011,
    72'b110000000000000000110000000000000000000000000000000000000000000000000000,
    72'b110000000000000111110000000000000000000000000000000000000000000000000000
};

const logic [0:8][0:3] ONE_BITMAP = {
    4'b0000,
    4'b1110,
    4'b0110,
    4'b0110,
    4'b0110,
    4'b0110,
    4'b1111,
    4'b0000,
    4'b0000
};

const logic [0:8][0:3] TWO_BITMAP = {
    4'b0000,
    4'b0110,
    4'b1001,
    4'b0011,
    4'b0110,
    4'b1100,
    4'b1111,
    4'b0000,
    4'b0000
};